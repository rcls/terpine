library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.defs.all;

entity cycle is
  generic (phase_init : natural range 0 to 3);
  port (R : out word_t;
        Din : in word_t;
        load : in std_logic;
        phase_advance : in std_logic;
        clk : in std_logic);
end cycle;

-- 'load' to 'A' is 6 cycle latency.
-- 'Din' to 'A' is 5 cycle latency.
-- 'phase_advance' to 'A' is 5 cycle latency.
-- Then 79 cycles to first result.
architecture cycle of cycle is
  function F0(B : word_t; C : word_t; D : word_t) return word_t is
  begin
      return (B and C) or (not B and D);
  end F0;

  function F1(B : word_t; C : word_t; D : word_t) return word_t is
  begin
      return B xor C xor D;
  end F1;

  function F2(B : word_t; C : word_t; D : word_t) return word_t is
  begin
      return (B and C) or (C and D) or (D and B);
  end F2;

  constant iA : word_t := x"67452301";
  constant iB : word_t := x"efcdab89";
  constant iC : word_t := x"98badcfe";
  constant iD : word_t := x"10325476";
  constant iE : word_t := x"c3d2e1f0";

  constant k0 : word_t := x"5a827999";
  constant k1 : word_t := x"6ed9eba1";
  constant k2 : word_t := x"8f1bbcdc";
  constant k3 : word_t := x"ca62c1d6";

  signal phase3 : natural range 0 to 3 := phase_init;
  signal munged_phase2 : natural range 0 to 3;

  signal A : word_t;
  signal C2 : word_t;
  signal D2 : word_t;
  signal I1 : word_t;
  signal I2 : word_t;
  signal I3 : word_t;

  signal init1_or_2 : boolean;
  signal init2_or_3 : boolean;
  --signal init3 : boolean;

  signal W : word_t;
  signal W2 : word_t;
  signal W3 : word_t;
  signal W8 : word_t;
  signal W14 : word_t;
  signal W15 : word_t;

  -- We split into 4 to rloc them seperately.
  signal W16a : unsigned(0 to 7);
  signal W16b : unsigned(0 to 7);
  signal W16c : unsigned(0 to 7);
  signal W16d : unsigned(0 to 7);

  signal pa : std_logic;
  signal ld : std_logic;

  attribute keep_hierarchy : string;
  attribute keep_hierarchy of cycle : architecture is "soft";

  attribute hu_set : string;
  attribute rloc : string;
  constant col8 : string :=
    "X1Y7 X1Y7 X1Y7 X1Y7 " &
    "X1Y6 X1Y6 X1Y6 X1Y6 " &
    "X1Y5 X1Y5 X1Y5 X1Y5 " &
    "X1Y4 X1Y4 X1Y4 X1Y4 " &
    "X1Y3 X1Y3 X1Y3 X1Y3 " &
    "X1Y2 X1Y2 X1Y2 X1Y2 " &
    "X1Y1 X1Y1 X1Y1 X1Y1 " &
    "X1Y0 X1Y0 X1Y0 X1Y0";
  attribute hu_set of I2 : signal is "I2_D2";
  attribute hu_set of D2 : signal is "I2_D2";
  attribute rloc of I2 : signal is col8;
  attribute rloc of D2 : signal is col8;

  attribute hu_set of A : signal is "A_W2";
  attribute hu_set of W2 : signal is "A_W2";
  attribute rloc of A : signal is col8;
  attribute rloc of W2 : signal is col8;

  attribute hu_set of W : signal is "W_W3";
  attribute hu_set of W3 : signal is "W_W3";
  attribute rloc of W : signal is col8;
  attribute rloc of W3 : signal is col8;

  attribute hu_set of I3 : signal is "I3_W15";
  attribute hu_set of W15 : signal is "I3_W15";
  attribute rloc of I3 : signal is col8;
  attribute rloc of W15 : signal is col8;

  attribute hu_set of W16a : signal is "W16a";
  attribute hu_set of W16b : signal is "W16b";
  attribute hu_set of W16c : signal is "W16c";
  attribute hu_set of W16d : signal is "W16d";
  attribute rloc of W16a : signal is "X0Y0";
  attribute rloc of W16b : signal is "X0Y0";
  attribute rloc of W16c : signal is "X0Y0";
  attribute rloc of W16d : signal is "X0Y0";

begin
  R <= A;

  d7_13 : entity work.double_delay generic map (7, 13)
    port map (w, w, w8, w14, clk);
  --d14_16 : entity work.double_delay generic map (13, 15)
  --  port map (w, w, w14, w16, clk);

  process
    variable kk : word_t;
    variable init1 : boolean;
    variable init2 : boolean;
    variable init3 : boolean;
  begin
    wait until rising_edge(clk);

    init1 := init1_or_2 and not init2_or_3;
    init2 := init1_or_2 and init2_or_3;
    init3 := init2_or_3 and not init1_or_2;

    -- 1 cycle latency into A.
    A <= (A rol 5) + I1;
    if init1 then
      A <= (iA rol 5) + F0(iB, iC, iD) - F0(iA, iB rol 30, iC) + I1;
    end if;

    -- 2 cycle latency into A.
    case munged_phase2 is -- 1 instead of 3; 3 means init1 or init2.
      when 0 => I1 <= F0(A, C2, D2) + I2;
      when 1 => I1 <= F1(A, C2, D2) + I2;
      when 2 => I1 <= F2(A, C2, D2) + I2;
      when 3 => I1 <= F0(iA, iB rol 30, iC) + I2;
    end case;

    -- Look aheads for these, and set up for init 1.
    C2 <= A rol 30;
    D2 <= C2;
    if init1 then
      C2 <= iA rol 30;
    end if;
    if init2 then
      C2 <= iB rol 30;
    end if;
    if init3 then
      C2 <= iC;
    end if;

    -- 3 cycle latency into A.
    I2 <= D2 + I3;
    if init3 then
      I2 <= iE + I3;
    end if;
    if init2 then
      I2 <= iD + I3;
    end if;

    if init2 or init3 then
      munged_phase2 <= 3;
    elsif phase3 = 3 then
      munged_phase2 <= 1;
    else
      munged_phase2 <= phase3;
    end if;

    -- 4 cycle latency into A.
    if pa = '1' then
      case phase3 is                    -- Look-ahead...
        when 0 => kk := k1;
        when 1 => kk := k2;
        when 2 => kk := k3;
        when 3 => kk := k0;
      end case;
    else
      case phase3 is
        when 0 => kk := k0;
        when 1 => kk := k1;
        when 2 => kk := k2;
        when 3 => kk := k3;
      end case;
    end if;
    I3 <= kk + W;

    if pa = '1' then
      if ld = '1' or phase3 = 3 then
        phase3 <= 0;
      else
        phase3 <= phase3 + 1;
      end if;
    end if;

    init2_or_3 <= (phase3 = 3 and pa = '1') or init3;
    init1_or_2 <= init2_or_3;

    -- 5 cycle latency into A.
    if ld = '1' then
      W <= Din;
    else
      W <= (W3 xor W8 xor W14 xor (W16d & W16c & W16b & W16a)) rol 1;
    end if;
    W2 <= W;
    W3 <= W2;
    W15 <= W14;
    W16d <= W15(31 downto 24);
    W16c <= W15(23 downto 16);
    W16b <= W15(15 downto  8);
    W16a <= W15( 7 downto  0);

    ld <= load;
    pa <= phase_advance;
  end process;
end cycle;
